/*
* Top level design of the FPGC6
*/
module FPGC6(
);


endmodule
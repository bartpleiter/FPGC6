/*
* B32P CPU
*/

module CPU(
    input clk, reset
);


endmodule
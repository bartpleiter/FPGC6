/*
* Timer
*/

module Timer(
    input clk, reset
);


endmodule
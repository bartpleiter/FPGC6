/*
* Instruction Decoder
*/

module InstructionDecoder(
    input clk, reset
);


endmodule
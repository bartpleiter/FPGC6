/*
* Stack
*/

module Stack (
    input clk, reset
);


endmodule
/*
* Control Unit
*/

module ControlUnit(
    input           clk, reset
);  


endmodule
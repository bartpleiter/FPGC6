/*
* ALU
*/

module ALU(
    input       [31:0]  a, b,
    input       [3:0]   opcode,
    output reg  [31:0]  y
);

endmodule
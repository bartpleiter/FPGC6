/*
* Register Bank
*/

module Regbank(
    input clk, reset
);


endmodule
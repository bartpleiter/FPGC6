/*
* L1 Cache
* Sits between Datamem or Instrmem and arbiter
*/
module L1cache(
);

endmodule